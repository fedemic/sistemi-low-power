A <= '1';
B <= '1';
S <= '1', '0' after 1 ns;
